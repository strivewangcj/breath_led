module led();



endmodule