module led(
input clk,
input rst_n


);



endmodule